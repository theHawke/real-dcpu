/**************************************************************************
 *  FPGA-implementation of the dcpu16
 *  Copyright (C) 2013  Hauke Neizel
 *
 *  This program is free software; you can redistribute it and/or modify
 *  it under the terms of the GNU General Public License as published by
 *  the Free Software Foundation; either version 2 of the License, or
 *  (at your option) any later version.
 *
 *  This program is distributed in the hope that it will be useful,
 *  but WITHOUT ANY WARRANTY; without even the implied warranty of
 *  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *  GNU General Public License for more details.
 *
 *  You should have received a copy of the GNU General Public License along
 *  with this program; if not, write to the Free Software Foundation, Inc.,
 *  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
 *
 */

module DEV_TEMPLATE (

	// CPU/Interrupt interactio ("Westbridge")
	
	
	// DMA ("Eastbridge")
	input DMA_CLOCK,
	input DMA_access, // whether this device has the access right this cycle
	output DMA_want, // whether this device needs DMA at the moment
	output [15:0] DMA_addr,
	output [15:0] DMA_out,
	output DMA_wren,
	input DMA_data

	// Device Specific I/O (clocks etc.)
	

);



endmodule

// modules for the direct memory access for devices
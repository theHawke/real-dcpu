// modules for the interrupt interaction between devices and the CPU